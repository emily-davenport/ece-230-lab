// Our top module is in our memory system because Vivado doesn't like me